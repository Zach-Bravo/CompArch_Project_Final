module RegDecoder (en,I,o);

input [4:0]I;
input en;

output reg [0:32] o;

//wire [4:0] W;
//assign I[4:0] = W[4:0];
//register_file (.I(I[4:0]));

		always @ (I or en) begin
			if (en==1'b1) begin
		
		 
				case (I)
			
					5'b00000 : o=32'b00000000000000000000000000000001;
					5'b00001 : o=32'b00000000000000000000000000000010;
					5'b00010 : o=32'b00000000000000000000000000000100;
					5'b00011 : o=32'b00000000000000000000000000001000;
					5'b00100 : o=32'b00000000000000000000000000010000;
					5'b00101 : o=32'b00000000000000000000000000100000;
					5'b00110 : o=32'b00000000000000000000000001000000;
					5'b00111 : o=32'b00000000000000000000000010000000;
					5'b01000 : o=32'b00000000000000000000000100000000;
					5'b01001 : o=32'b00000000000000000000001000000000;
					5'b01010 : o=32'b00000000000000000000010000000000;
					5'b01011 : o=32'b00000000000000000000100000000000;
					5'b01100 : o=32'b00000000000000000001000000000000;
					5'b01101 : o=32'b00000000000000000010000000000000;
					5'b01110 : o=32'b00000000000000000100000000000000;
					5'b01111 : o=32'b00000000000000001000000000000000;
					5'b10000 : o=32'b00000000000000010000000000000000;
					5'b10001 : o=32'b00000000000000100000000000000000;
					5'b10010 : o=32'b00000000000001000000000000000000;
					5'b10011 : o=32'b00000000000010000000000000000000;
					5'b10100 : o=32'b00000000000100000000000000000000;
					5'b10101 : o=32'b00000000001000000000000000000000;
					5'b10110 : o=32'b00000000010000000000000000000000;
					5'b10111 : o=32'b00000000100000000000000000000000;
					5'b11000 : o=32'b00000001000000000000000000000000;
					5'b11001 : o=32'b00000010000000000000000000000000;
					5'b11010 : o=32'b00000100000000000000000000000000;
					5'b11011 : o=32'b00001000000000000000000000000000;
					5'b11100 : o=32'b00010000000000000000000000000000;
					5'b11101 : o=32'b00100000000000000000000000000000;
					5'b11110 : o=32'b01000000000000000000000000000000;
					5'b11111 : o=32'b10000000000000000000000000000000;
					default : o=32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

	endcase	 
		end
			end

endmodule 	

/*module decoder2to4(in, o);
input [1:0] in;
output reg [3:0] o;

always @ (in)begin
	case(in)
		2'b00 : o= 4'b0001;
		2'b01 : o= 4'b0010;
		2'b10 : o= 4'b0100;
		2'b11 : o= 4'b1000;	
default : o = 4'bxxxx;
	
endcase
end 		
endmodule*/